module Controller (
);
    
endmodule